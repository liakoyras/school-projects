library verilog;
use verilog.vl_types.all;
entity keyboard_tb is
end keyboard_tb;
